[Grass]
id=grass
textureFilename=grass_0.png

[Water]
id=water
textureFilename=water_0.png

[Swamp]
id=swamp
textureFilename=blob.png
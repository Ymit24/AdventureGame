[Grassland]
id=grassland_basic
textureFilename=grassland_bullet.png
projectileBehavior=straight
projectileEmitter=single
firingRate=1.25
damage=

[Spider]
id=spider_attack
textureFilename=bullet_0.png
projectileBehavior=sine
projectileEmitter=triple
firingRate=.6
damage=5

[PurpleWand]
id=purple_wand
textureFilename=bullet_0.png
projectileBehavior=straight
projectileEmitter=single
firingRate=0.25
damage=1

[GreenStaff]
id=green_staff
textureFilename=bullet_1.png
projectileBehavior=sine
projectileEmitter=double_together
firingRate=0.45
damage=3

[BlueWand]
id=blue_wand
textureFilename=bullet_2.png
projectileBehavior=straight
projectileEmitter=triple
firingRate=1
damage=6

[YellowStaff]
id=yellow_staff
textureFilename=bullet_2.png
projectileBehavior=sine
projectileEmitter=circle
firingRate=0.6
damage=13
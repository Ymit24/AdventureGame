[BlobEasy]
id=blob_easy
moveSpeed=0.45
health=6
textureFilename=blob_0.png
xpDrop=1
weaponId=grassland_basic

[BlobMedium]
id=blob_med
moveSpeed=0.55
health=44
textureFilename=blob_1.png
xpDrop=3
weaponId=grassland_basic

[BlobHard]
id=blob_hard
moveSpeed=0.65
health=123
textureFilename=blob_2.png
xpDrop=9
weaponId=grassland_basic

[ImpersonatorEasy]
id=impersonator_easy
moveSpeed=2.25
health=8
textureFilename=impersonator_0.png
xpDrop=2
weaponId=grassland_basic

[ImpersonatorMedium]
id=impersonator_med
moveSpeed=3
health=64
textureFilename=impersonator_1.png
xpDrop=6
weaponId=grassland_basic

[ImpersonatorHard]
id=impersonator_hard
moveSpeed=3.4
health=154
textureFilename=impersonator_2.png
xpDrop=13
weaponId=grassland_basic

[Spider]
id=spider
moveSpeed=2.5
health=425
textureFilename=swamp/spider.png
xpDrop=27
weaponId=grassland_basic

[SwampBlob]
id=swamp_blob
moveSpeed=2
health=640
textureFilename=swamp/swamp_blob.png
xpDrop=40
weaponId=grassland_basic
[Grass]
id=grass
textureFilename=sprites/grass_0.png

[Water]
id=water
textureFilename=sprites/water_0.png

[Swamp]
id=swamp
textureFilename=sprites/blob.png
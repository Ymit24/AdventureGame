[SimpleWand]
id=simple_wand
textureFilename=bullet_0.png
projectileBehavior=straight
projectileEmitter=single
firingRate=0.25
damage=1

[SpecialStaff]
id=spec_staff
textureFilename=bullet_1.png
projectileBehavior=sine
projectileEmitter=double_together
firingRate=0.45
damage=3

[Thing]
id=some_weapon
textureFilename=bullet_2.png
projectileBehavior=straight
projectileEmitter=triple
firingRate=1
damage=6
[Tree]
id=tree
name=Grassland Tree
textureFilename=tree_0.png
collision=true
[BlobEasy]
id=blob_easy
moveSpeed=0.45
health=6
textureFilename=blob_0.png
xpDrop=1

[BlobMedium]
id=blob_med
moveSpeed=0.55
health=44
textureFilename=blob_1.png
xpDrop=3

[BlobHard]
id=blob_hard
moveSpeed=0.65
health=123
textureFilename=blob_2.png
xpDrop=9

[ImpersonatorEasy]
id=impersonator_easy
moveSpeed=2.25
health=8
textureFilename=impersonator_0.png
xpDrop=2

[ImpersonatorMedium]
id=impersonator_med
moveSpeed=3
health=64
textureFilename=impersonator_1.png
xpDrop=6

[ImpersonatorHard]
id=impersonator_hard
moveSpeed=3.4
health=154
textureFilename=impersonator_2.png
xpDrop=13
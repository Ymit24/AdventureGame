[Grass]
id=grass
textureFilename=grass_0.png

[Water]
id=water
textureFilename=water_0.png

[Path]
id=path
textureFilename=path_0.png
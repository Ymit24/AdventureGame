[Grass]
id=grass
textureFilename=grass_0.png
isWalkable=true

[Water]
id=water
textureFilename=water_0.png
isWalkable=false

[Path]
id=path
textureFilename=path_0.png
isWalkable=true

[Swamp]
id=swamp
textureFilename=swamp/swamp_0.png
isWalkable=true
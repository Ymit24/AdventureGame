[Grassland]
id=grassland_basic
textureFilename=grassland_bullet.png
projectileBehavior=straight
projectileEmitter=single
firingRate=1.25
damage=2

[MidLand]
id=midland_basic
textureFilename=bullet_2.png
projectileBehavior=straight
projectileEmitter=double
firingRate=0.75
damage=4

[MidLandAlt]
id=midland_alt
textureFilename=bullet_1.png
projectileBehavior=straight
projectileEmitter=circle
firingRate=0.5
damage=3

[Highland]
id=highland_basic
textureFilename=bullet_2.png
projectileBehavior=sine
projectileEmitter=double_together
firingRate=0.3
damage=4

[Highland]
id=highland_alt
textureFilename=bullet_1.png
projectileBehavior=straight
projectileEmitter=triple
firingRate=0.25
damage=3

[Spider]
id=spider_attack
textureFilename=bullet_0.png
projectileBehavior=sine
projectileEmitter=triple
firingRate=.6
damage=5

[PurpleWand]
id=purple_wand
textureFilename=bullet_0.png
projectileBehavior=straight
projectileEmitter=single
firingRate=0.45
damage=2

[BlueWand]
id=blue_wand
textureFilename=bullet_2.png
projectileBehavior=straight
projectileEmitter=triple
firingRate=.6
damage=6

[GreenStaff]
id=green_staff
textureFilename=bullet_1.png
projectileBehavior=sine
projectileEmitter=double_together
firingRate=0.17
damage=13

[YellowStaff]
id=yellow_staff
textureFilename=bullet_2.png
projectileBehavior=sine
projectileEmitter=circle
firingRate=0.25
damage=25